module hello;
  initial 
    begin
      $display("Verilog is Hardware Description Language. Hello! World.");
      $finish ;
    end
endmodule
